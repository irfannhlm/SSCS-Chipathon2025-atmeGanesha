* Testbench
.param fnoicor = 0
.param sw_stat_mismatch = 0
.lib "/foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice" typical
.include "ptl_mux.spice"  *Include spice netlist

* Drives power supply
VDD VDD 0 3.3V

* Drives input signal
VINS S 0 PULSE(0 3.3 0n 0.1n 0.1n 5n 10n)
VINA A 0 PULSE(0 3.3 0n 0.1n 0.1n 10n 20n)
VINB B 0 PULSE(0 3.3 0n 0.1n 0.1n 20n 40n) 

* Transient analysis
.tran 1n 50n
.option TEMP=25

.control
  run
  plot v(S)+10.5 v(A)+7.0 v(B)+3.5 v(OUT)
.endc

.end

